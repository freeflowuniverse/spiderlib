module spider