module auth

[noinit]
struct AuthServer {

}



pub fn new() {}