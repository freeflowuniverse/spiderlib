module vapi

struct APIConfig {
	
}

struct API {

}