module partials

struct List {
}
