module ssg

// fn gen
