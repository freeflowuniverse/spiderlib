module session