module main 

// fn (app PaymentApp) fulfill_ourphone_order(session Session) {
// 	//todo: implement
// }