module spider

fn install_tailwind() {

}

fn load_tailwind() {

}

fn preprocess_tailwind() {

}