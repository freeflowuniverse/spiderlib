module tailwindui
