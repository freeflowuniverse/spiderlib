module main

import 