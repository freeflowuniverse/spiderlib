module ssg


// pub fn build(path string) {
// 	new


// }

