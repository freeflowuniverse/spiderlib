module ssg

// fn gen