module uikit2
