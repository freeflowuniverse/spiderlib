module flowbite

