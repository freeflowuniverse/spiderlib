module main

// import vweb

// pub struct TailwindUI {
// 	vweb.Context
// }
