module tailwindui

import freeflowuniverse.spiderlib.uikit

struct Page {
	uikit.Page
}