module tailwindui