module uikitweb

// import vweb

// pub struct TailwindUI {
// 	vweb.Context
// }
