module partials

pub struct Table {
pub:
	headers []string
	rows [][]string
}