module uikit2