module ssg

fn parse_content() {
}
