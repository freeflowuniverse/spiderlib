module vapi


// generates api key
fn generate_key() {
	
}

// verifies api key
fn verify_key() bool {
	return true
}