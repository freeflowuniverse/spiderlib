module stripeclient

pub fn (client StripeClient) get_customer(customer_id string) Customer {
	return Customer{}
}