module uikit