module dependency

