module server

pub fn (mut app App) refresh() vweb.Result {
}
