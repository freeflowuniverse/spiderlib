module main

struct Registrar {
    registrations map[string]Registration
}

struct Registration {
    name string
    email string
}

pub fn (mut model Registrar) register(name string, email string) {
    model.registrations << 
}

pub fn (model Registrar) get_registrations(name string, email string) {

}