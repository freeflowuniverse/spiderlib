module api

struct APIConfig {
}

struct API {
}
