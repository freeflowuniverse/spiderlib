module main

// import
