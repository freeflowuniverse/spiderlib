module partials

struct List {
	
}